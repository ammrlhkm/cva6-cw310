`define BERGEN
// include KINTEX7 specific code (relevant for KC705, GENESYSII,...)
`define ARIANE_DATA_WIDTH 64

// Instantiate protocl checker
// `define PROTOCOL_CHECKER
